//
// File : ppi_tx_if.svh
//
// Created:
//          by HDL Designers Team
//          of Electronics Design Center "OhT"
//          www.overhitech.com
//
//
// File Description:
//
//% Интерфейс CSi (bidirectional)
//

`ifndef __CSI_BIDIR_IF_SVH__
    `define __CSI_BIDIR_IF_SVH__

`include "vivo_env_structural_defines.svh"
    
    //----------------------------------------------------------------------------------------------------------------------
    // CSI PPI-bidir interface
    //----------------------------------------------------------------------------------------------------------------------

interface oht_vivo_csi_bidir_if#(int LANE_N = `OHT_VIVO_CSI_LANES_MAX);

    //------------------------------------------------------------------------------------------------------------------
    // Pin declaration
    //------------------------------------------------------------------------------------------------------------------
    
    wire clk_n;
    wire clk_p;
    wire [LANE_N-1:0] data_n;
    wire [LANE_N-1:0] data_p;

    //------------------------------------------------------------------------------------------------------------------
    // Test wires
    //------------------------------------------------------------------------------------------------------------------
    
    //------------------------------------------------------------------------------------------------------------------
    // Modports
    //------------------------------------------------------------------------------------------------------------------
    
    modport checker_mp (
        input clk_n,
        input clk_p,
        input data_n,
        input data_p
    );
    
endinterface

`endif // __CSI_BIDIR_IF_SVH__